library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package dmem is
    type data_out is array(0 to 479) of std_logic_vector(7 downto 0);
end package;

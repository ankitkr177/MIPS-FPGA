library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package IMem is
    type instr_out is array(0 to 651) of std_logic_vector(7 downto 0);
end package;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.std_logic_unsigned.all;
USE IEEE.STD_LOGIC_ARITH.ALL;
use work.IMem.all;

entity InstructionMemory is
    Port ( PC : in STD_LOGIC_VECTOR (31 downto 0);
           Instr : inout STD_LOGIC_VECTOR (31 downto 0));
end InstructionMemory;

architecture Behavioral of InstructionMemory is

constant IMem1 : instr_out := instr_out'(
"00110000","00000000","00000000","10010011", -- JUMPS TO INSTRUCTION 147PLACEHOLDER FOR JUMP
"00011100","00011111","00000000","00100000", --lw $0, $31, 32   // load $31 with (1000...000) from dmem(32)
"00000100","00001010","00000000","00011010", --addi $0, $10, 26  //$10 stores value 26  changed
"00000100","00001011","00000000","00000100", --addi $0, $11, 4   //$11 stores value 4   changed
"00000100","00001100","00000000","01001110", --addi $0, $12, 78  //$12 stores value 78
"00011100","11000011","00000000","00000000", --lw $6, $3, 0      //load S(0) to $3
"00000000","01100001","01001000","00000001", --add $3, $1, $9    //$9=A+S(0)
"00000001","00100010","01001000","00000001", --add $9, $2, $9    //$9=A+B+S(0)
"00000001","00111111","11110000","00000101", --*and $9, $31, $30 (1000...00) -- take the first digit in r30
"00010101","00101001","00000000","00000001", --shl $9, $9, 1     //$9=(A+B+skey(0))<<<1 
"00101000","00011110","00000000","00000001", --*beq $30, $0, 1 (subi $8, $8, 1 )      // Check if r31 has msb 1 or 0
"00000101","00101001","00000000","00000001", --*addi $9, $9, 1      // if msb 1 add 1 to shifted value
"00000001","00111111","11110000","00000101", --*and $9, $31, $30 (1000...00) -- take the first digit in r30
"00010101","00101001","00000000","00000001", --shl $9, $9, 1     //$9=(A+B+skey(0))<<<1 
"00101000","00011110","00000000","00000001", --*beq $30, $0, 1 (subi $8, $8, 1 )      // Check if r31 has msb 1 or 0
"00000101","00101001","00000000","00000001", --*addi $9, $9, 1      // if msb 1 add 1 to shifted value
"00000001","00111111","11110000","00000101", --*and $9, $31, $30 (1000...00) -- take the first digit in r30
"00010101","00101001","00000000","00000001", --shl $9, $9, 1     //$9=(A+B+skey(0))<<<1 
"00101000","00011110","00000000","00000001", --*beq $30, $0, 1 (subi $8, $8, 1 )      // Check if r31 has msb 1 or 0
"00000101","00101001","00000000","00000001", --*addi $9, $9, 1      // if msb 1 add 1 to shifted value
"00000000","00001001","00001000","00000001", --add $0, $9, $1    //put A value back to $1
"00100000","11000001","00000000","00000000", --sw $6, $1, 0      //store the A value back to S(0)
"00000000","00100010","01000000","00000001", --add $1, $2, $8    //$8=A+B
"00001101","00001000","00000000","00011111", --andi $8, $8, 31   //put last five bits of A+B into $8
"00011100","11100100","00000000","00011010", --lw $7, $4, 26     //$4=ukey(0)
"00000000","10000001","01001000","00000001", --add $4, $1, $9    //$9=A+ukey(0)
"00000001","00100010","01001000","00000001", --add $9, $2, $9    //$9=A+B+ukey(0)
"00101000","00001000","00000000","00000110", --beq $0, $8, 6 (add $0, $9, $2 )    //check whether $9 has finished shift 
"00000001","00111111","11110000","00000101", --*and $9, $31, $30 (1000...00) -- take the first digit in r30
"00010101","00101001","00000000","00000001", --shl $9, $9, 1     //$9=(A+B+ukey(0))<<<1
"00101000","00011110","00000000","00000001", --*beq $30, $0, 1 (subi $8, $8, 1 )      // Check if r31 has msb 1 or 0
"00000101","00101001","00000000","00000001", --*addi $9, $9, 1      // if msb 1 add 1 to shifted value
"00001001","00001000","00000000","00000001", --subi $8, $8, 1    
"00101100","00001000","00000000","00001100", --bne $0, $8, 12 (jump intgr 14)    //check whether $9 has finished shift, if not go back to shift ////changed
"00000000","00001001","00010000","00000001", --add $0, $9, $2    //put B value back to $2
"00100000","11100010","00000000","00011010", --sw $7, $2, 26     //store B value back to ukey(0)
"00000100","11000110","00000000","00000001", --addi $6, $6, 1    //$6 is i counter  changed
"00000100","11100111","00000000","00000001", --addi $7, $7, 1    //$7 is j counter  changed
"00101100","11001010","00000000","00000001", --bne $6, $10, 1 (bne $7, $11, 1)    //check i counter
"00000000","11000110","00110000","00000011", --sub $6, $6, $6    //if i counter is 26, set back to 0
"00101100","11101011","00000000","00000001", --bne $7, $11, 1  (addi $5, $5, 1)   //check j counter
"00000000","11100111","00111000","00000011", --sub $7, $7, $7    //if j counter is 4, set back to 0
"00000100","10100101","00000000","00000001", --addi $5, $5, 1    //$5 is counter for key expansion
"00101100","10101100","00000000","00000001", --bne $5, $12, 1 (jump top) //if $5 is not 78, go back to do the loop
"00110000","00000000","00000000","10011010", --halt REPLACED WITH JUMP 47 (sub $5, $5, $5) to encryption
"00110000","00000000","00000000","00000101", --jump top 5 (lw $6, $3, 0)
"00110000","00000000","00000000","00011011", -- jump intgr 27 (beq $0, $8, 6)
"00000000","10100101","00101000","00000011", --*sub $5, $5, $5  -----ENCRYPTION  
"00000000","11000110","00110000","00000011", --*sub $6, $6, $6  
"00000000","11100111","00111000","00000011", --*sub $7, $7, $7   
"00000001","10001100","01100000","00000011", --*sub $12, $12, $12  
"00011100","00000001","00000000","00011110", --*lw $0, $1, 30       //$1=A
"00011100","00000010","00000000","00011111", --*lw $0, $2, 31       //$2=B
"00011100","00011111","00000000","00100000", --*lw $0, $31, 32   // load $31 with (1000...000) from dmem(32)
"00011100","00000011","00000000","00000000", --lw $0, $3, 0       //$3=S(0)
"00011100","00000100","00000000","00000001", --lw $0, $4, 1       //$4=S(1)
"00000000","00100011","00001000","00000001", --add $1, $3, $1     //$1=A+S(0)
"00000000","01000100","00010000","00000001", --add $2, $4, $2     //$2=B+S(1)
"00000100","00001100","00000000","00001100", --addi $0, $12, 12   //store value 12 in $12
"00000000","00100010","00100000","00000111", --or $1, $2, $4      //$4=A or B
"00000000","00100010","00101000","00000101", --and $1, $2, $5     //$5=A and B
"00000000","10000101","00100000","00000011", --sub $4, $5, $4     //$4=(A or B)-(A and B)=A xor B
"00001100","01000101","00000000","00011111", --andi $2, $5, 31    //put the last five bits of B into $5
"00000100","11000110","00000000","00000001", --addi $6, $6, 1     //$6 is the i counter
"00101000","00000101","00000000","00000110", --beq $0, $5, 6 (SHL $6, $7, 1)     //check wether shift has finished ---check it
"00000000","10011111","11110000","00000101", --*and $4, $31, $30 (1000...00) -- take the first digit in r30
"00010100","10000100","00000000","00000001", --SHL $4, $4, 1      //if not, $4=(A xor B)<<<1
"00101000","00011110","00000000","00000001", --*beq $30, $0, 1 (subi $8, $8, 1 )      // Check if r31 has msb 1 or 0
"00000100","10000100","00000000","00000001", --*addi $4, $4, 1      // if msb 1 add 1 to shifted value
"00001000","10100101","00000000","00000001", --SUBI $5, $5, 1 
"00101100","00000101","00000000","00010101", --BNE $0, $5, 21 (jmp 17)    //check wether shift has finished ----check it
"00010100","11000111","00000000","00000001", --SHL $6, $7, 1      //$7=$6*2
"00011100","11100011","00000000","00000000", --LW $7, $3, 0       //$3=S(2)
"00000000","10000011","00001000","00000001", --ADD $4, $3, $1     //$1=a_rot+S(2), put A value back to $1
"00000000","00100010","00100000","00000111", --OR $1, $2, $4      //$4=A or B
"00000000","00100010","00101000","00000101", --and $1, $2, $5     //$5=A and B
"00000000","10000101","00100000","00000011", --sub $4, $5, $4     //$4=(A or B)-(A and B)=A xor B
"00001100","00100101","00000000","00011111", --andi $1, $5, 31    //put the last five bits of A into $5
"00101000","00000101","00000000","00000110", --beq $0, $5, 6 (addi $7, $7, 1)     //check wether shift has finished
"00000000","10011111","11110000","00000101", --*and $4, $31, $30 (1000...00) -- take the first digit in r30
"00010100","10000100","00000000","00000001", --shl $4, $4, 1      //if not, $4=(A xor B)<<<1
"00101000","00011110","00000000","00000001", --*beq $30, $0, 1 (subi $8, $8, 1 )      // Check if r31 has msb 1 or 0
"00000100","10000100","00000000","00000001", --*addi $4, $4, 1      // if msb 1 add 1 to shifted value
"00001000","10100101","00000000","00000001", --subi $5, $5, 1
"00101100","00000101","00000000","00001000", --bne $0, $5, 8  (jmp 31)   //check wether shift has finished
"00000100","11100111","00000000","00000001", --addi $7, $7, 1     //$7=2*i+1
"00011100","11100011","00000000","00000000", --lw $7, $3, 0       //$3=S(3)
"00000000","10000011","00010000","00000001", --add $4, $3, $2     //$2=A+B, put B value back to $2
"00101101","10000110","00000000","00000101", --bne $12, $6, 5 (jmp 5)  //check if the 12 loop has finished, if not go back
"00100000","00000001","00000000","00100001", --sw $0, $1, 33      //store A value into data memory
"00100000","00000010","00000000","00100010", --sw $0, $2, 34      //store B value into data memory
"00110000","00000000","00000000","10011101", --hal REPLACED WITH JMP FAILSAFE
"00110000","00000000","00000000","01000000", --jmp 64 (beq $0, $5, 6 upper )
"00110000","00000000","00000000","01001110", --jmp 78 (beq $0, $5, 6 lower)
"00110000","00000000","00000000","00111011", --jmp 59 (or $1, $2, $4 )
"00000001","10001100","01100000","00000011", --*sub $12, $12, $12 ------DECRYPTION
"00000011","10111101","11101000","00000011", --*sub $29, $29, $29  
"00000100","00011101","00000000","00100000", --*addi $0, $29, 32 
"00011100","00000001","00000000","00100001", --*lw $0, $1, 33       //$1=A
"00011100","00000010","00000000","00100010", --*lw $0, $2, 34       //$2=B
"00011100","00011111","00000000","00100000", --*lw $0, $31, 32   // load $31 with (1000...000) from dmem(32)
"00000100","00001100","00000000","00001100", --addi $0, $12, 12   //store value 12 into $12, i_counter
"00010101","10001101","00000000","00000001", --shl $12, $13, 1    //$13=2*i
"00000101","10101110","00000000","00000001", --addi $13, $14, 1   //$14=2*i+1 
"00011101","11000011","00000000","00000000", --lw $14, $3, 0      //$3=S(25)
"00000000","01000011","00010000","00000011", --sub $2, $3, $2     //$2=B-S(25)
"00001100","00100100","00000000","00011111", --andi $1, $4, 31    //put the last five bits of A into $4
"00000011","10100100","00100000","00000011", --*sub $29, $4, $4 
"00101011","10100100","00000000","00000110", --beq $29, $4, 6 (or $1, $2, $5 )  //check if the loop has finished
"00000000","01011111","11110000","00000101", --*and $2, $31, $30 (1000...00) -- take the first digit in r30
"00010100","01000010","00000000","00000001", --shl $2, $2, 1      //if not, $2=(B-S(25))>>>1
"00101000","00011110","00000000","00000001", --*beq $30, $0, 1 (subi $4, $4, 1 ) // Check if r31 has msb 1 or 0
"00000100","01000010","00000000","00000001", --*addi $2, $2, 1      // if msb 1 add 1 to shifted value
"00001000","10000100","00000000","00000001", --subi $4, $4, 1
"00101100","00000100","00000000","00011101", --bne $0, $4, 29 (jmp 13)    //check if the loop has finished
"00000000","00100010","00101000","00000111", --or $1, $2, $5      //$5=((B-S(25))>>>A) or A
"00000000","00100010","00110000","00000101", --and $1, $2, $6     //$6=((B-S(25))>>>A) and A
"00000000","10100110","00010000","00000011", --sub $5, $6, $2     //$2=((B-S(25))>>>A) xor A
"00000000","01100011","00011000","00000011", --sub $3, $3, $3     //clear $3
"00011101","10100011","00000000","00000000", --lw $13, $3, 0      //$3=S(24)
"00000000","00100011","00001000","00000011", --sub $1, $3, $1     //$1=A-S(24)
"00001100","01000100","00000000","00011111", --andi $2, $4, 31    //put the last five bits of B into $4
"00000011","10100100","00100000","00000011", --*sub $29, $4, $4 
"00101011","10100100","00000000","00000110", --beq $29, $4, 6 (or $1, $2, $5)  //check if the loop has finished
"00000000","00111111","11110000","00000101", --*and $1, $31, $30 (1000...00) -- take the first digit in r30
"00010100","00100001","00000000","00000001", --shl $1, $1, 1      //if not, $1=(A-S(24))>>>1
"00101000","00011110","00000000","00000001", --*beq $30, $0, 1 (subi $4, $4, 1 ) // Check if r31 has msb 1 or 0
"00000100","00100001","00000000","00000001", --*addi $1, $1, 1      // if msb 1 add 1 to shifted value
"00001000","10000100","00000000","00000001", --subi $4, $4, 1
"00101100","00000100","00000000","00001111", --bne $0, $4, 15 (jmp 28)  //check if the loop has finished
"00000000","00100010","00101000","00000111", --or $1, $2, $5      //$5=((A-S(24))>>>B) or B
"00000000","00100010","00110000","00000101", --and $1, $2, $6     //$6=((A-S(24))>>>B) and B
"00000000","10100110","00001000","00000011", --sub $5, $6, $1     //$6=((A-S(24))>>>B) xor B
"00001001","10001100","00000000","00000001", --subi $12, $12, 1   //reduce 1 from i counter
"00101101","10000000","00000000","00001011", --bne $12, $0, 11 (jmp 7)   //check if 12 loop has finished, if not, go back to loop
"00000000","01100011","00011000","00000011", --sub $3, $3, $3     //if yes, clear $3
"00011100","00000011","00000000","00000001", --lw $0, $3, 1       //$3=S(1)
"00000000","01000011","00010000","00000011", --sub $2, $3, $2     //$2=B-S(1)
"00000000","01100011","00011000","00000011", --sub $3, $3, $3
"00011100","00000011","00000000","00000000", --lw $0, $3, 0       //$3=S(0)
"00000000","00100011","00001000","00000011", --sub $1, $3, $1     //$1=A-S(0)
"00100000","00000001","00000000","00100011", --*******sw $0, $1, 35      //store A value to data memory
"00100000","00000010","00000000","00100100", --*******sw $0, $2, 36      //store B value to data memory
"00110000","00000000","00000000","10100000", --hal REPLACED WITH JUMP
"00110000","00000000","00000000","01101100", --jmp 108 (beq $29, $4, 6 upper)
"00110000","00000000","00000000","01111011", --jmp 123 (beq $29, $4, 6 lower)
"00110000","00000000","00000000","01100110", --jmp 102 (shl $12, $13, 1)  
"00101100","00010000","00000000","00000011", --**bne $0, $16, 3 
"00101100","00010001","00000000","00000011", --**bne $0, $17, 3
"00101100","00010010","00000000","00000011", --**bne $0, $18, 3  
"00110000","00000000","00000000","10010011", --**jmp instr 147
"00110000","00000000","00000000","00000001", --**jmp to key expansion
"00110000","00000000","00000000","00101111", --**jmp to encryption
"00110000","00000000","00000000","01011111", --**jmp to decryption
"00101100","00010000","00000000","00000001", --**bne $16, $0, 1 ---jumps here after key expansion (FAILSAFE)
"00110000","00000000","00000000","10010011", --**jmp instr 147
"00110000","00000000","00000000","10011010", --**jmp 154loop failsafe for key expansion until $16 is set to approriate 
"00101100","00010001","00000000","00000001", --**bne $17, $0, 1 ---jumps here after encryption (FAILSAFE)
"00110000","00000000","00000000","10010011", --**jmp instr 147
"00110000","00000000","00000000","10011101", --**jmp 157 loop failsafe for encryption until $17 is set to approriate 
"00101100","00010010","00000000","00000001", --**bne $18, $0, 1 ---jumps here after decryption (FAILSAFE)
"00110000","00000000","00000000","10010011", --**jmp instr 147
"00110000","00000000","00000000","10100000"); --**jmp 160 loop failsafe for dencryption until $18 is set to approriate 
 

--constant IMem1 : instr_out := instr_out'(
--"00110000","00000000","00000000","00000001", -- PLACEHOLDER FOR JUMP
--"00011100","00011111","00000000","00100000", --lw $0, $31, 32   // load $31 with (1000...000) from dmem(32)
--"00000100","00001010","00000000","00011010", --addi $0, $10, 26  //$10 stores value 26  changed
--"00000100","00001011","00000000","00000100", --addi $0, $11, 4   //$11 stores value 4   changed
--"00000100","00001100","00000000","01001110", --addi $0, $12, 78  //$12 stores value 78
--"00011100","11000011","00000000","00000000", --lw $6, $3, 0      //load S(0) to $3
--"00000000","01100001","01001000","00000001", --add $3, $1, $9    //$9=A+S(0)
--"00000001","00100010","01001000","00000001", --add $9, $2, $9    //$9=A+B+S(0)
--"00000001","00111111","11110000","00000101", --*and $9, $31, $30 (1000...00) -- take the first digit in r30
--"00010101","00101001","00000000","00000001", --shl $9, $9, 1     //$9=(A+B+skey(0))<<<1 
--"00101000","00011110","00000000","00000001", --*beq $30, $0, 1 (subi $8, $8, 1 )      // Check if r31 has msb 1 or 0
--"00000101","00101001","00000000","00000001", --*addi $9, $9, 1      // if msb 1 add 1 to shifted value
--"00000001","00111111","11110000","00000101", --*and $9, $31, $30 (1000...00) -- take the first digit in r30
--"00010101","00101001","00000000","00000001", --shl $9, $9, 1     //$9=(A+B+skey(0))<<<1 
--"00101000","00011110","00000000","00000001", --*beq $30, $0, 1 (subi $8, $8, 1 )      // Check if r31 has msb 1 or 0
--"00000101","00101001","00000000","00000001", --*addi $9, $9, 1      // if msb 1 add 1 to shifted value
--"00000001","00111111","11110000","00000101", --*and $9, $31, $30 (1000...00) -- take the first digit in r30
--"00010101","00101001","00000000","00000001", --shl $9, $9, 1     //$9=(A+B+skey(0))<<<1 
--"00101000","00011110","00000000","00000001", --*beq $30, $0, 1 (subi $8, $8, 1 )      // Check if r31 has msb 1 or 0
--"00000101","00101001","00000000","00000001", --*addi $9, $9, 1      // if msb 1 add 1 to shifted value
--"00000000","00001001","00001000","00000001", --add $0, $9, $1    //put A value back to $1
--"00100000","11000001","00000000","00000000", --sw $6, $1, 0      //store the A value back to S(0)
--"00000000","00100010","01000000","00000001", --add $1, $2, $8    //$8=A+B
--"00001101","00001000","00000000","00011111", --andi $8, $8, 31   //put last five bits of A+B into $8
--"00011100","11100100","00000000","00011010", --lw $7, $4, 26     //$4=ukey(0)
--"00000000","10000001","01001000","00000001", --add $4, $1, $9    //$9=A+ukey(0)
--"00000001","00100010","01001000","00000001", --add $9, $2, $9    //$9=A+B+ukey(0)
--"00101000","00001000","00000000","00000110", --beq $0, $8, 6 (add $0, $9, $2 )    //check whether $9 has finished shift 
--"00000001","00111111","11110000","00000101", --*and $9, $31, $30 (1000...00) -- take the first digit in r30
--"00010101","00101001","00000000","00000001", --shl $9, $9, 1     //$9=(A+B+ukey(0))<<<1
--"00101000","00011110","00000000","00000001", --*beq $30, $0, 1 (subi $8, $8, 1 )      // Check if r31 has msb 1 or 0
--"00000101","00101001","00000000","00000001", --*addi $9, $9, 1      // if msb 1 add 1 to shifted value
--"00001001","00001000","00000000","00000001", --subi $8, $8, 1    
--"00101100","00001000","00000000","00001100", --bne $0, $8, 12 (jump intgr 14)    //check whether $9 has finished shift, if not go back to shift ////changed
--"00000000","00001001","00010000","00000001", --add $0, $9, $2    //put B value back to $2
--"00100000","11100010","00000000","00011010", --sw $7, $2, 26     //store B value back to ukey(0)
--"00000100","11000110","00000000","00000001", --addi $6, $6, 1    //$6 is i counter  changed
--"00000100","11100111","00000000","00000001", --addi $7, $7, 1    //$7 is j counter  changed
--"00101100","11001010","00000000","00000001", --bne $6, $10, 1 (bne $7, $11, 1)    //check i counter
--"00000000","11000110","00110000","00000011", --sub $6, $6, $6    //if i counter is 26, set back to 0
--"00101100","11101011","00000000","00000001", --bne $7, $11, 1  (addi $5, $5, 1)   //check j counter
--"00000000","11100111","00111000","00000011", --sub $7, $7, $7    //if j counter is 4, set back to 0
--"00000100","10100101","00000000","00000001", --addi $5, $5, 1    //$5 is counter for key expansion
--"00101100","10101100","00000000","00000001", --bne $5, $12, 1 (jump top) //if $5 is not 78, go back to do the loop
--"00110000","00000000","00000000","00101111", --halt REPLACED WITH JUMP 47 (sub $5, $5, $5) to encryption
--"00110000","00000000","00000000","00000101", --jump top 5 (lw $6, $3, 0)
--"00110000","00000000","00000000","00011011", -- jump intgr 27 (beq $0, $8, 6)begin
--"00000000","10100101","00101000","00000011", --*sub $5, $5, $5  -----ENCRYPTION  
--"00000000","11000110","00110000","00000011", --*sub $6, $6, $6  
--"00000000","11100111","00111000","00000011", --*sub $7, $7, $7   
--"00000001","10001100","01100000","00000011", --*sub $12, $12, $12  
--"00011100","00000001","00000000","00011110", --*lw $0, $1, 30       //$1=A
--"00011100","00000010","00000000","00011111", --*lw $0, $2, 31       //$2=B
--"00011100","00011111","00000000","00100000", --*lw $0, $31, 32   // load $31 with (1000...000) from dmem(32)
--"00011100","00000011","00000000","00000000", --lw $0, $3, 0       //$3=S(0)
--"00011100","00000100","00000000","00000001", --lw $0, $4, 1       //$4=S(1)
--"00000000","00100011","00001000","00000001", --add $1, $3, $1     //$1=A+S(0)
--"00000000","01000100","00010000","00000001", --add $2, $4, $2     //$2=B+S(1)
--"00000100","00001100","00000000","00001100", --addi $0, $12, 12   //store value 12 in $12
--"00000000","00100010","00100000","00000111", --or $1, $2, $4      //$4=A or B
--"00000000","00100010","00101000","00000101", --and $1, $2, $5     //$5=A and B
--"00000000","10000101","00100000","00000011", --sub $4, $5, $4     //$4=(A or B)-(A and B)=A xor B
--"00001100","01000101","00000000","00011111", --andi $2, $5, 31    //put the last five bits of B into $5
--"00000100","11000110","00000000","00000001", --addi $6, $6, 1     //$6 is the i counter
--"00101000","00000101","00000000","00000110", --beq $0, $5, 6 (SHL $6, $7, 1)     //check wether shift has finished ---check it
--"00000000","10011111","11110000","00000101", --*and $4, $31, $30 (1000...00) -- take the first digit in r30
--"00010100","10000100","00000000","00000001", --SHL $4, $4, 1      //if not, $4=(A xor B)<<<1
--"00101000","00011110","00000000","00000001", --*beq $30, $0, 1 (subi $8, $8, 1 )      // Check if r31 has msb 1 or 0
--"00000100","10000100","00000000","00000001", --*addi $4, $4, 1      // if msb 1 add 1 to shifted value
--"00001000","10100101","00000000","00000001", --SUBI $5, $5, 1 
--"00101100","00000101","00000000","00010101", --BNE $0, $5, 21 (jmp 17)    //check wether shift has finished ----check it
--"00010100","11000111","00000000","00000001", --SHL $6, $7, 1      //$7=$6*2
--"00011100","11100011","00000000","00000000", --LW $7, $3, 0       //$3=S(2)
--"00000000","10000011","00001000","00000001", --ADD $4, $3, $1     //$1=a_rot+S(2), put A value back to $1
--"00000000","00100010","00100000","00000111", --OR $1, $2, $4      //$4=A or B
--"00000000","00100010","00101000","00000101", --and $1, $2, $5     //$5=A and B
--"00000000","10000101","00100000","00000011", --sub $4, $5, $4     //$4=(A or B)-(A and B)=A xor B
--"00001100","00100101","00000000","00011111", --andi $1, $5, 31    //put the last five bits of A into $5
--"00101000","00000101","00000000","00000110", --beq $0, $5, 6 (addi $7, $7, 1)     //check wether shift has finished
--"00000000","10011111","11110000","00000101", --*and $4, $31, $30 (1000...00) -- take the first digit in r30
--"00010100","10000100","00000000","00000001", --shl $4, $4, 1      //if not, $4=(A xor B)<<<1
--"00101000","00011110","00000000","00000001", --*beq $30, $0, 1 (subi $8, $8, 1 )      // Check if r31 has msb 1 or 0
--"00000100","10000100","00000000","00000001", --*addi $4, $4, 1      // if msb 1 add 1 to shifted value
--"00001000","10100101","00000000","00000001", --subi $5, $5, 1
--"00101100","00000101","00000000","00001000", --bne $0, $5, 8  (jmp 31)   //check wether shift has finished
--"00000100","11100111","00000000","00000001", --addi $7, $7, 1     //$7=2*i+1
--"00011100","11100011","00000000","00000000", --lw $7, $3, 0       //$3=S(3)
--"00000000","10000011","00010000","00000001", --add $4, $3, $2     //$2=A+B, put B value back to $2
--"00101101","10000110","00000000","00000101", --bne $12, $6, 5 (jmp 5)  //check if the 12 loop has finished, if not go back
--"00100000","00000001","00000000","00011110", --sw $0, $1, 30      //store A value into data memory
--"00100000","00000010","00000000","00011111", --sw $0, $2, 31      //store B value into data memory
--"11111100","00000000","00000000","00000000", --hal
--"00110000","00000000","00000000","01000000", --jmp 64 (beq $0, $5, 6 upper )
--"00110000","00000000","00000000","01001110", --jmp 78 (beq $0, $5, 6 lower)
--"00110000","00000000","00000000","00111011"); --jmp 59 (or $1, $2, $4 )

begin

Instr <= (IMem1(conv_integer(unsigned(PC)))) &  (IMem1(conv_integer(unsigned(PC+1)))) &
         (IMem1(conv_integer(unsigned(PC+2)))) &  (IMem1(conv_integer(unsigned(PC+3))));

end Behavioral;
